-- FIFOWRAPPER.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FIFOWRAPPER is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity FIFOWRAPPER;

architecture rtl of FIFOWRAPPER is
	component FIFOWRAPPER_FIFO_WRAPPER_0 is
	end component FIFOWRAPPER_FIFO_WRAPPER_0;

begin

	fifo_wrapper_0 : component FIFOWRAPPER_FIFO_WRAPPER_0
		port map (
		);

end architecture rtl; -- of FIFOWRAPPER
