----------------------------------------------------------------------------------
--
-- Company:          Flat Earth, Inc.
-- Author/Engineer:	Ross K. Snider
--
-- Create Date:      09/09/2016
--
-- Design Name:      AD1939.vhd  
--       				
-- Description:      The AD1939 component does the following:
--									1. Initializes all the AD1939 registers (Configure AD1939_init.mif to set hard coded power up register settings.  This can be generated by the Matlab file AD1939_init.m)
--									2. Allows individual register writes (to change volume, sample rate, etc.)
--                         3. Provids a simple data interface for reading & writing CODEC data
--                         4. AD1939 is configured in 24-bit normal stereo serial mode (see page 15 of AD1939 data sheet)
--
-- Target Device(s): Altera DE0-Nano-Soc Evaluation Board
-- Tool versions:    Quartus Prime 16.0
--
-- Dependencies:     AD1939.vhd
--                       AD1939_Control.vhd
--                       AD1939_Data.vhd
--
-- Revisions:        1.0 (File Created)
--
-- Additional Comments: 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity AD1939 is
	port
	(	
		AD1939_SPI_CLK : in  std_logic; -- SPI Clock that must be < 10 MHz
		reset          : in  std_logic; -- system reset
		AD1939_MCLK    : out std_logic; -- 12.8 MHz Master Clock from AD1939 crystal
		state_monitor  : out std_logic_vector (3 downto 0);  -- debug
		----------------------------------------------------------------------------------------------------------------
		-- Physical Layer : signals to SPI port
		-- Signals to/from AD1939 SPI Control Port (data direction from AD1939 perspective), connection to physical pins on AD1939
		-- 10 MHz CCLK max (see page 7 of AD1939 data sheet)
		-- CIN data is 24-bits (see page 14 of AD1939 data sheet)
		-- CLATCH_n must have pull-up resistor so that AD1939 recognizes presence of SPI controller on power-up
		----------------------------------------------------------------------------------------------------------------
		AD1939_SPI_CIN      : out std_logic;  		 -- SPI Control Data Input to AD1939 pin 30 CIN
		AD1939_SPI_COUT     : in  std_logic;       -- SPI Control Data output from AD1939 pin 31 COUT
		AD1939_SPI_CCLK     : out std_logic;       -- SPI Control Clock Input to AD1939 pin 34 CCLK
		AD1939_SPI_CLATCH_n : out std_logic;       -- SPI Latch for control data, input to AD1939 pin 35 CLATCH_n (active low)
		-------------------------------------------------------------------------------------------------------------------------------------
		-- Physical Layer : signals to serial data port on AD1939
		-- Signals to/from AD1939 Serial Data Port (from ADCs/to DACs), i.e. connection to physical pins on AD1939
		-------------------------------------------------------------------------------------------------------------------------------------
		AD1939_ADC_SDATA1          : in     std_logic;   -- Serial data from AD1939 pin 27 ASDATA1, ADC1 24-bit normal stereo serial mode
		AD1939_ADC_SDATA2          : in     std_logic;   -- Serial data from AD1939 pin 26 ASDATA2, ADC2 24-bit normal stereo serial mode
		AD1939_ADC_BCLK            : in     std_logic;   -- Serial data from AD1939 pin 28 ABCLK, Bit Clock for ADCs (Master Mode)
		AD1939_ADC_LRCLK           : in     std_logic;   -- Serial data from AD1939 pin 29 ALRCLK, LR Clock for ADCs (Master Mode)
		--
		AD1939_DAC_SDATA1          : out    std_logic;   -- Serial data to AD1939 pin 20 DSDATA1, DAC1 24-bit normal stereo serial mode
		AD1939_DAC_SDATA2          : out    std_logic;   -- Serial data to AD1939 pin 19 DSDATA2, DAC2 24-bit normal stereo serial mode
		AD1939_DAC_SDATA3          : out    std_logic;   -- Serial data to AD1939 pin 18 DSDATA3, DAC3 24-bit normal stereo serial mode
		AD1939_DAC_SDATA4          : out    std_logic;   -- Serial data to AD1939 pin 15 DSDATA4, DAC4 24-bit normal stereo serial mode
		AD1939_DAC_BCLK            : out    std_logic;   -- Serial data to AD1939 pin 21 DBCLK, Bit Clock for DACs (Slave Mode)
		AD1939_DAC_LRCLK           : out    std_logic;   -- Serial data to AD1939 pin 22 DLRCLK, LR Clock for DACs (Slave Mode)
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- Abstracted register interface to AD1939
		-- Simple interface to read/write AD1939 register data
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		AD1939_Reg_Addr				: in 		std_logic_vector (4 downto 0);   -- Address of AD1939 Register to be read/written (there are 17 registers)
		AD1939_Reg_Write_Data		: in 		std_logic_vector (7 downto 0);   -- Data to be written to AD1939 Register
		AD1939_Reg_Write_Start  	: in 		std_logic;                       -- Initiates the register write when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data			: out		std_logic_vector (7 downto 0);   -- Data read from AD1939 Register
		AD1939_Reg_Read_Start	   : in 		std_logic;                       -- Initiates the register read when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data_Ready	: out		std_logic;   							-- Clock pulse signifies data read from AD1939 Register and is ready to be captured
		AD1939_Reg_Busy	         : out 	std_logic;                       -- read or write is occurring, any new read/write will be ignored 
		-----------------------------------------------------------------------------------------------------------
		-- Abstracted data channels, i.e. interface to data plane 
		-- Interface for reading and writing AD1939 ADC/DAC (sample) 24-bit data (data is in 2's complement form)???
		-----------------------------------------------------------------------------------------------------------
		-- Data from ADCs
		AD1939_Data_ADC1_Left   : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC1_Right  : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC2_Left   : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC2_Right  : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADCs_ready  : out std_logic;                        -- pulse 1 BCLK period wide signifies data is ready to read from ADCs (this pulse occurs at the sample rate Fs) 	
      --	Data to DACs	
		AD1939_Data_DAC1_Left   : in std_logic_vector (23 downto 0);    -- On the rising edge of the DAC_LRCLK, these DAC signals will be captured 
		AD1939_Data_DAC1_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC2_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC2_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC3_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC3_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC4_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC4_Right  : in std_logic_vector (23 downto 0)
	);
end AD1939;

architecture behavioral of AD1939 is
	
	----------------------------------------------------------------------------------------------------------
	-- AD1939_control
	-- Component that initializes the AD1939 register settings and allows individual register read/writes.
	----------------------------------------------------------------------------------------------------------
	component AD1939_control 
		port (
		AD1939_SPI_CLK : in  std_logic; -- SPI Clock (also component clock) that must be <= 10 MHz
		reset          : in  std_logic; -- system reset
		state_monitor  : out std_logic_vector (3 downto 0);  -- debug
		----------------------------------------------------------------------------------------------------------------
		-- Signals to/from AD1939 SPI Control Port (data direction from AD1939 perspective)
		-- 10 MHz CCLK max (see page 7 of AD1939 data sheet)
		-- CIN data is 24-bits (see page 14 of AD1939 data sheet)
		-- CLATCH_n must have pull-up resistor so that AD1939 recognizes presence of SPI controller on power-up
		----------------------------------------------------------------------------------------------------------------
		AD1939_SPI_CIN      : out std_logic;  		 -- SPI Control Data Input to AD1939 pin 30 CIN
		AD1939_SPI_COUT     : in  std_logic;       -- SPI Control Data output from AD1939 pin 31 COUT
		AD1939_SPI_CCLK     : out std_logic;       -- SPI Control Clock Input to AD1939 pin 34 CCLK
		AD1939_SPI_CLATCH_n : out std_logic;       -- SPI Latch for control data, input to AD1939 pin 35 CLATCH_n (active low)
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- Simple interface to read/write AD1939 register data
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		AD1939_Reg_Addr				: in 		std_logic_vector (4 downto 0);   -- Address of AD1939 Register to be read/written (there are 17 registers)
		AD1939_Reg_Write_Data		: in 		std_logic_vector (7 downto 0);   -- Data to be written to AD1939 Register
		AD1939_Reg_Write_Start  	: in 		std_logic;                       -- Initiates the register write when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data			: out		std_logic_vector (7 downto 0);   -- Data read from AD1939 Register
		AD1939_Reg_Read_Start	   : in 		std_logic;                       -- Initiates the register read when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data_Ready	: out		std_logic;   							-- Clock pulse signifies data read from AD1939 Register and is ready to be captured
		AD1939_Reg_Busy	         : out 	std_logic                        -- read or write is occurring, any new read/write will be ignored 
		 );
	end component;
	
	----------------------------------------------------------------------------------------------------------
	-- AD1939_data
	-- Component that converts the ADC serial data into parallel and parallel DAC data to serial
	----------------------------------------------------------------------------------------------------------
	component AD1939_data is
		port
		(	
			reset          : in  std_logic; -- system reset
			AD1939_MCLK    : out std_logic; -- 12.8 MHz Master Clock from AD1939 crystal
			-------------------------------------------------------------------------------------------------------------------------------------
			-- Physical Layer : signals to serial data port on AD1939
			-- Signals to/from AD1939 Serial Data Port (from ADCs/to DACs), i.e. connection to physical pins on AD1939
			-------------------------------------------------------------------------------------------------------------------------------------
			AD1939_ADC_SDATA1          : in     std_logic;   -- Serial data from AD1939 pin 27 ASDATA1, ADC1 24-bit normal stereo serial mode
			AD1939_ADC_SDATA2          : in     std_logic;   -- Serial data from AD1939 pin 26 ASDATA2, ADC2 24-bit normal stereo serial mode
			AD1939_ADC_BCLK            : in     std_logic;   -- Serial data from AD1939 pin 28 ABCLK, Bit Clock for ADCs (Master Mode)
			AD1939_ADC_LRCLK           : in     std_logic;   -- Serial data from AD1939 pin 29 ALRCLK, LR Clock for ADCs (Master Mode)
			--
			AD1939_DAC_SDATA1          : out    std_logic;   -- Serial data to AD1939 pin 20 DSDATA1, DAC1 24-bit normal stereo serial mode
			AD1939_DAC_SDATA2          : out    std_logic;   -- Serial data to AD1939 pin 19 DSDATA2, DAC2 24-bit normal stereo serial mode
			AD1939_DAC_SDATA3          : out    std_logic;   -- Serial data to AD1939 pin 18 DSDATA3, DAC3 24-bit normal stereo serial mode
			AD1939_DAC_SDATA4          : out    std_logic;   -- Serial data to AD1939 pin 15 DSDATA4, DAC4 24-bit normal stereo serial mode
			AD1939_DAC_BCLK            : out    std_logic;   -- Serial data to AD1939 pin 21 DBCLK, Bit Clock for DACs (Slave Mode)
			AD1939_DAC_LRCLK           : out    std_logic;   -- Serial data to AD1939 pin 22 DLRCLK, LR Clock for DACs (Slave Mode)
			-----------------------------------------------------------------------------------------------------------
			-- Abstracted data channels, i.e. interface to FPGA data plane 
			-- Interface for reading and writing AD1939 ADC/DAC (sample) 24-bit data (data is in 2's complement form)???
			-----------------------------------------------------------------------------------------------------------
			-- Data from ADCs
			AD1939_Data_ADC1_Left   : out std_logic_vector(23 downto 0); 
			AD1939_Data_ADC1_Right  : out std_logic_vector(23 downto 0); 
			AD1939_Data_ADC2_Left   : out std_logic_vector(23 downto 0); 
			AD1939_Data_ADC2_Right  : out std_logic_vector(23 downto 0); 
			AD1939_Data_ADCs_ready  : out std_logic;                        -- pulse 1 BCLK period wide signifies data is ready to read from ADCs (this pulse occurs at the sample rate Fs) 	
			--	Data to DACs	
			AD1939_Data_DAC1_Left   : in std_logic_vector(23 downto 0);    -- On the rising edge of the DAC_LRCLK, these DAC signals will be captured 
			AD1939_Data_DAC1_Right  : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC2_Left   : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC2_Right  : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC3_Left   : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC3_Right  : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC4_Left   : in std_logic_vector(23 downto 0); 
			AD1939_Data_DAC4_Right  : in std_logic_vector(23 downto 0)
		);
	end component;
				
begin

	--------------------------------------------------------------------------------------
	-- Component that controls AD1939
	--------------------------------------------------------------------------------------
	u1 : AD1939_control
	port map (
		AD1939_SPI_CLK => AD1939_SPI_CLK, -- SPI Clock (also component clock) that must be <= 10 MHz
		reset          => reset,          -- system reset
		state_monitor  => state_monitor, -- debug
		----------------------------------------------------------------------------------------------------------------
		-- Exported signals to/from AD1939 SPI Control Port (data direction from AD1939 perspective)
		-- 10 MHz CCLK max (see page 7 of AD1939 data sheet)
		-- CIN data is 24-bits (see page 14 of AD1939 data sheet)
		-- CLATCH_n must have pull-up resistor so that AD1939 recognizes presence of SPI controller on power-up
		----------------------------------------------------------------------------------------------------------------
		AD1939_SPI_CIN      =>  AD1939_spi_CIN,		 -- SPI Control Data Input to AD1939 pin 30 CIN
		AD1939_SPI_COUT     =>  AD1939_spi_COUT,     -- SPI Control Data output from AD1939 pin 31 COUT
		AD1939_SPI_CCLK     =>  AD1939_spi_CCLK,     -- SPI Control Clock Input to AD1939 pin 34 CCLK
		AD1939_SPI_CLATCH_n =>  AD1939_spi_CLATCH_n,     -- SPI Latch for control data, input to AD1939 pin 35 CLATCH_n (active low)
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- Simple interface to read/write AD1939 register data
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		AD1939_Reg_Addr					=> AD1939_Reg_Addr, -- Address of AD1939 Register to be read/written (there are 17 registers)
		AD1939_Reg_Write_Data			=> AD1939_Reg_Write_Data, -- Data to be written to AD1939 Register
		AD1939_Reg_Write_Start  		=> AD1939_Reg_Write_Start,                     -- Initiates the register write when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data				=> AD1939_Reg_Read_Data, -- Data read from AD1939 Register
		AD1939_Reg_Read_Start			=> AD1939_Reg_Read_Start,                   -- Initiates the register read when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data_Ready		=> AD1939_Reg_Read_Data_Ready, 							-- Clock pulse signifies data read from AD1939 Register and is ready to be captured
		AD1939_Reg_Busy	      		=> AD1939_Reg_Busy                     -- read or write is occurring, any new read/write will be ignored 
	 );
	
	
	----------------------------------------------------------------------------------------------------------
	-- AD1939_data
	-- Component that converts the ADC serial data into parallel and parallel DAC data to serial
	----------------------------------------------------------------------------------------------------------
	u2 : AD1939_data
	port map (
		reset          => reset, -- system reset
		AD1939_MCLK    => AD1939_MCLK, -- 12.8 MHz Master Clock from AD1939 crystal
		-------------------------------------------------------------------------------------------------------------------------------------
		-- Physical Layer : signals to serial data port on AD1939
		-- Signals to/from AD1939 Serial Data Port (from ADCs/to DACs), i.e. connection to physical pins on AD1939
		-------------------------------------------------------------------------------------------------------------------------------------
		AD1939_ADC_SDATA1          => AD1939_ADC_SDATA1,   -- Serial data from AD1939 pin 27 ASDATA1, ADC1 24-bit normal stereo serial mode
		AD1939_ADC_SDATA2          => AD1939_ADC_SDATA2,   -- Serial data from AD1939 pin 26 ASDATA2, ADC2 24-bit normal stereo serial mode
		AD1939_ADC_BCLK            => AD1939_ADC_BCLK,   -- Serial data from AD1939 pin 28 ABCLK, Bit Clock for ADCs (Master Mode)
		AD1939_ADC_LRCLK           => AD1939_ADC_LRCLK,   -- Serial data from AD1939 pin 29 ALRCLK, LR Clock for ADCs (Master Mode)
		--
		AD1939_DAC_SDATA1          => AD1939_DAC_SDATA1,  -- Serial data to AD1939 pin 20 DSDATA1, DAC1 24-bit normal stereo serial mode
		AD1939_DAC_SDATA2          => AD1939_DAC_SDATA2,  -- Serial data to AD1939 pin 19 DSDATA2, DAC2 24-bit normal stereo serial mode
		AD1939_DAC_SDATA3          => AD1939_DAC_SDATA3,  -- Serial data to AD1939 pin 18 DSDATA3, DAC3 24-bit normal stereo serial mode
		AD1939_DAC_SDATA4          => AD1939_DAC_SDATA4,  -- Serial data to AD1939 pin 15 DSDATA4, DAC4 24-bit normal stereo serial mode
		AD1939_DAC_BCLK            => AD1939_DAC_BCLK,  -- Serial data to AD1939 pin 21 DBCLK, Bit Clock for DACs (Slave Mode)
		AD1939_DAC_LRCLK           => AD1939_DAC_LRCLK,  -- Serial data to AD1939 pin 22 DLRCLK, LR Clock for DACs (Slave Mode)
		-----------------------------------------------------------------------------------------------------------
		-- Abstracted data channels, i.e. interface to FPGA data plane 
		-- Interface for reading and writing AD1939 ADC/DAC (sample) 24-bit data (data is in 2's complement form)???
		-----------------------------------------------------------------------------------------------------------
		-- Data from ADCs
		AD1939_Data_ADC1_Left   => AD1939_Data_ADC1_Left,
		AD1939_Data_ADC1_Right  => AD1939_Data_ADC1_Right,
		AD1939_Data_ADC2_Left   => AD1939_Data_ADC2_Left,
		AD1939_Data_ADC2_Right  => AD1939_Data_ADC2_Right,
		AD1939_Data_ADCs_ready  => AD1939_Data_ADCs_ready,                       -- pulse 1 BCLK period wide signifies data is ready to read from ADCs (this pulse occurs at the sample rate Fs) 	
		--	Data to DACs	
		AD1939_Data_DAC1_Left   => AD1939_Data_DAC1_Left,   -- On the rising edge of the DAC_LRCLK, these DAC signals will be captured 
		AD1939_Data_DAC1_Right  => AD1939_Data_DAC1_Right,
		AD1939_Data_DAC2_Left   => AD1939_Data_DAC2_Left,
		AD1939_Data_DAC2_Right  => AD1939_Data_DAC2_Right,
		AD1939_Data_DAC3_Left   => AD1939_Data_DAC3_Left,
		AD1939_Data_DAC3_Right  => AD1939_Data_DAC3_Right,
		AD1939_Data_DAC4_Left   => AD1939_Data_DAC4_Left,
		AD1939_Data_DAC4_Right  => AD1939_Data_DAC4_Right
	);
		
end behavioral;
	
	
	
	
	
	
	