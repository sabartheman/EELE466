----------------------------------------------------------------------------------
--
-- Company:          Flat Earth, Inc.
-- Author/Engineer:	Ross K. Snider
--
-- Create Date:      09/09/2016
--
-- Design Name:      AD1939_top.vhd  
--       				
-- Description:      The AD1939_top component does the following:
--									1. Initializes all the AD1939 registers (Configure AD1939_init.mif to set hard coded power up register settings.  This can be generated by the Matlab file AD1939_init.m)
--									2. Allows individual register writes (to change volume, sample rate, etc.)
--                         3. Provids a simple data interface for reading & writing CODEC data
--                         4. AD1939 is configured in 24-bit normal stereo serial mode (see page 15 of AD1939 data sheet)
--
-- Target Device(s): Altera DE0-Nano-Soc Evaluation Board
-- Tool versions:    Quartus Prime 16.0
--
-- Dependencies:     AD1939_top.vhd
--                       AD1939_Control.vhd
--                       AD1939_Data.vhd
--
-- Revisions:        1.0 (File Created)
--
-- Additional Comments: 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity AD1939_top is
	port
	(	
		clk			   : in  std_logic; -- system clock
		reset          : in  std_logic; -- system reset
		AD1939_MCLK    : out std_logic; -- 12.8 MHz Master Clock from AD1939 crystal
		AD1939_SPI_CLK : in  std_logic; -- SPI Clock that must be < 10 MHz
		AD1939_RST_n   : in  std_logic; -- AD1939 Power Down Reset (Active Low) to AD1939 pin 14 PD_n/RST_n 
		AD1939_pin_14  : out std_logic;
		----------------------------------------------------------------------------------------------------------------
		-- Signals to/from AD1939 SPI Control Port (data direction from AD1939 perspective)
		-- 10 MHz CCLK max (see page 7 of AD1939 data sheet)
		-- CIN data is 24-bits (see page 14 of AD1939 data sheet)
		-- CLATCH_n must have pull-up resistor so that AD1939 recognizes presence of SPI controller on power-up
		----------------------------------------------------------------------------------------------------------------
		AD1939_SPI_CIN      : out std_logic;  		 -- SPI Control Data Input to AD1939 pin 30 CIN
		AD1939_SPI_COUT     : in  std_logic;       -- SPI Control Data output from AD1939 pin 31 COUT
		AD1939_SPI_CCLK     : out std_logic;       -- SPI Control Clock Input to AD1939 pin 34 CCLK
		AD1939_SPI_CLATCH_n : out std_logic;       -- SPI Latch for control data, input to AD1939 pin 35 CLATCH_n (active low)
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- Simple interface to read/write AD1939 register data
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		AD1939_Reg_Addr				: in 		std_logic_vector (4 downto 0);   -- Address of AD1939 Register to be read/written (there are 17 registers)
		AD1939_Reg_Write_Data		: in 		std_logic_vector (7 downto 0);   -- Data to be written to AD1939 Register
		AD1939_Reg_Write_Start  	: in 		std_logic;                       -- Initiates the register write when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data			: out		std_logic_vector (7 downto 0);   -- Data read from AD1939 Register
		AD1939_Reg_Read_Start	   : in 		std_logic;                       -- Initiates the register read when asserted, must be deasserted to return from busy
		AD1939_Reg_Busy	         : out 	std_logic;                       -- read or write is occurring, any new read/write will be ignored 
		-------------------------------------------------------------------------------------------------------------------------------------
		-- Signals to/from AD1939 Serial Data Port (from ADCs/to DACs)
		-------------------------------------------------------------------------------------------------------------------------------------
		AD1939_ADC_SDATA1          : in     std_logic;   -- Serial data from AD1939 pin 27 ASDATA1, ADC1 24-bit normal stereo serial mode
		AD1939_ADC_SDATA2          : in     std_logic;   -- Serial data from AD1939 pin 26 ASDATA2, ADC2 24-bit normal stereo serial mode
		AD1939_ADC_BCLK            : in     std_logic;   -- Serial data from AD1939 pin 28 ABCLK, Bit Clock for ADCs (Master Mode)
		AD1939_ADC_LRCLK           : in     std_logic;   -- Serial data from AD1939 pin 29 ALRCLK, LR Clock for ADCs (Master Mode)
		--
		AD1939_DAC_SDATA1          : out    std_logic;   -- Serial data to AD1939 pin 20 DSDATA1, DAC1 24-bit normal stereo serial mode
		AD1939_DAC_SDATA2          : out    std_logic;   -- Serial data to AD1939 pin 19 DSDATA2, DAC2 24-bit normal stereo serial mode
		AD1939_DAC_SDATA3          : out    std_logic;   -- Serial data to AD1939 pin 18 DSDATA3, DAC3 24-bit normal stereo serial mode
		AD1939_DAC_SDATA4          : out    std_logic;   -- Serial data to AD1939 pin 15 DSDATA4, DAC4 24-bit normal stereo serial mode
		AD1939_DAC_BCLK            : out    std_logic;   -- Serial data to AD1939 pin 21 DBCLK, Bit Clock for DACs (Slave Mode)
		AD1939_DAC_LRCLK           : out    std_logic;   -- Serial data to AD1939 pin 22 DLRCLK, LR Clock for DACs (Slave Mode)
		-----------------------------------------------------------------------------------------------------------
		-- Interface for reading and writing AD1939 ADC/DAC (sample) 24-bit data (data is in 2's complement form)???
		-----------------------------------------------------------------------------------------------------------
		AD1939_Data_ADC1_Left   : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC1_Right  : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC2_Left   : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADC2_Right  : out std_logic_vector (23 downto 0); 
		AD1939_Data_ADCs_ready  : out std_logic;                        -- pulse 1 BCLK period wide signifies data is ready to read from ADCs (this pulse occurs at the sample rate Fs) 	
      --		
		AD1939_Data_DAC1_Left   : in std_logic_vector (23 downto 0);    -- On the rising edge of the DAC_LRCLK, these DAC signals will be captured 
		AD1939_Data_DAC1_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC2_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC2_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC3_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC3_Right  : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC4_Left   : in std_logic_vector (23 downto 0); 
		AD1939_Data_DAC5_Right  : in std_logic_vector (23 downto 0)
	);
end AD1939_top;

architecture behavioral of AD1939_top is
	
	----------------------------------------------------------------------------------------------------------
	-- AD1939_control
	-- Component that initializes the AD1939 register settings and allows individual register read/writes.
	----------------------------------------------------------------------------------------------------------
	component AD1939_control 
		port (
		clk			   : in  std_logic; -- system clock
		reset          : in  std_logic; -- system reset
		AD1939_SPI_CLK : in  std_logic; -- SPI Clock that must be < 10 MHz
		AD1939_RST_n   : in std_logic;  -- AD1939 Power Down Reset (Active Low) to AD1939 pin 14 PD_n/RST_n 
		AD1939_pin_14  : out std_logic;
		----------------------------------------------------------------------------------------------------------------
		-- Signals to/from AD1939 SPI Control Port (data direction from AD1939 perspective)
		-- 10 MHz CCLK max (see page 7 of AD1939 data sheet)
		-- CIN data is 24-bits (see page 14 of AD1939 data sheet)
		-- CLATCH_n must have pull-up resistor so that AD1939 recognizes presence of SPI controller on power-up
		----------------------------------------------------------------------------------------------------------------
		AD1939_SPI_CIN      : out std_logic;  		 -- SPI Control Data Input to AD1939 pin 30 CIN
		AD1939_SPI_COUT     : in  std_logic;       -- SPI Control Data output from AD1939 pin 31 COUT
		AD1939_SPI_CCLK     : out std_logic;       -- SPI Control Clock Input to AD1939 pin 34 CCLK
		AD1939_SPI_CLATCH_n : out std_logic;       -- SPI Latch for control data, input to AD1939 pin 35 CLATCH_n (active low)
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- Simple interface to read/write AD1939 register data
		----------------------------------------------------------------------------------------------------------------------------------------------------------------
		AD1939_Reg_Addr				: in 		std_logic_vector (4 downto 0);   -- Address of AD1939 Register to be read/written (there are 17 registers)
		AD1939_Reg_Write_Data		: in 		std_logic_vector (7 downto 0);   -- Data to be written to AD1939 Register
		AD1939_Reg_Write_Start  	: in 		std_logic;                       -- Initiates the register write when asserted, must be deasserted to return from busy
		AD1939_Reg_Read_Data			: out		std_logic_vector (7 downto 0);   -- Data read from AD1939 Register
		AD1939_Reg_Read_Start	   : in 		std_logic;                       -- Initiates the register read when asserted, must be deasserted to return from busy
		AD1939_Reg_Busy	         : out 	std_logic                        -- read or write is occurring, any new read/write will be ignored 
		 );
	end component;
	
--	component WM8731_Data 
--		port (
--				clk		: 	in 	std_logic;  -- DE2 board system 50 MHz clock 
--				reset 	: 	in		std_logic;  -- DE2 system reset				
--				-- WM8731 serial data signals
--				BCLK	 	: 	in 	std_logic;  -- Bit Clock coming from WM8731 (Master Mode - See figure 30 p. 37 of WM8731 datasheet) 
--				ADCLRC 	:  in 	std_logic;  -- Pulse 1 BCLK wide signifying start of data (DSP Mode - See figure 29 p. 34 of WM8731 datasheet)
--				ADCDAT 	: 	in		std_logic;  -- Serial data from ADC (Bit length assumed to be 24 bits, bit length set in IWL in register 7, see table on p. 50 of datasheet) 
--				DACLRC 	:  in 	std_logic;  -- Pulse 1 BCLK wide signifying start of data capture (DSP Mode - See figure 29 p. 34 of WM8731 datasheet)
--				DACDAT 	: 	out	std_logic;  -- Serial data to DAC (Bit length assumed to be 24 bits, bit length set in IWL in register 7, see table on p. 50 of datasheet) 
--				-- Data from ADC (in 2's complement form)
--				WM8731_Data_from_ADC_Left  : out std_logic_vector (23 downto 0); 
--				WM8731_Data_from_ADC_Right : out std_logic_vector (23 downto 0); 
--				WM8731_Data_from_ADC_ready : out std_logic; -- pulse 1 BCLK period wide signifying data is ready to read (this pulse occurs at the sample rate, i.e. Fs) 				
--				-- Data to DAC (in 2's complement form)
--				WM8731_Data_to_DAC_Left  : in std_logic_vector (23 downto 0); -- On the rising edge of the DACLRC Pulse, these output registers will be captured into an internal register and send out DACDAT
--				WM8731_Data_to_DAC_Right : in std_logic_vector (23 downto 0)
--		 );
--	end component;
				
begin

	--------------------------------------------------------------------------------------
	-- Component that controls AD1939
	--------------------------------------------------------------------------------------
	u1: AD1939_control 
	port map (
		clk			   			=> clk,
		reset          			=> reset, 
		AD1939_SPI_CLK 			=> AD1939_SPI_CLK,
		AD1939_RST_n   			=> AD1939_RST_n,
		AD1939_pin_14  			=> AD1939_pin_14,
		AD1939_SPI_CIN      		=> AD1939_SPI_CIN,
		AD1939_SPI_COUT     		=> AD1939_SPI_COUT,
		AD1939_SPI_CCLK     		=> AD1939_SPI_CCLK,
		AD1939_SPI_CLATCH_n 		=> AD1939_SPI_CLATCH_n,
		AD1939_Reg_Addr			=> AD1939_Reg_Addr,
		AD1939_Reg_Write_Data	=> AD1939_Reg_Write_Data,
		AD1939_Reg_Write_Start  => AD1939_Reg_Write_Start,
		AD1939_Reg_Read_Data		=> AD1939_Reg_Read_Data,
		AD1939_Reg_Read_Start	=> AD1939_Reg_Read_Start,
		AD1939_Reg_Busy	      => AD1939_Reg_Busy
    );
	
--	u3: WM8731_Data 
--	port map(
--			clk								=> MCLK,
--			reset 							=> reset,
--			BCLK	 							=> BCLK,
--			ADCLRC 							=> ADCLRC,
--			ADCDAT 							=> ADCDAT,
--			DACLRC 							=> DACLRC,
--			DACDAT 							=> DACDAT,
--			WM8731_Data_from_ADC_Left  => WM8731_Data_from_ADC_Left,
--			WM8731_Data_from_ADC_Right => WM8731_Data_from_ADC_Right,
--			WM8731_Data_from_ADC_ready => WM8731_Data_from_ADC_ready,
--			WM8731_Data_to_DAC_Left  	=> WM8731_Data_to_DAC_Left,
--			WM8731_Data_to_DAC_Right 	=> WM8731_Data_to_DAC_Right
--	);
		
end behavioral;
	
	
	
	
	
	
	