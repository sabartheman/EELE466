-- fifo_wrapper.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fifo_wrapper is
	port (
		clk_clk                                      : in  std_logic                     := '0';             --                        clk.clk
		fifo_wrapper_0_conduit_end_writebyteenable_n : in  std_logic_vector(3 downto 0)  := (others => '0'); -- fifo_wrapper_0_conduit_end.writebyteenable_n
		fifo_wrapper_0_conduit_end_readdata          : out std_logic_vector(3 downto 0);                     --                           .readdata
		fifo_wrapper_0_s1_address                    : in  std_logic_vector(4 downto 0)  := (others => '0'); --          fifo_wrapper_0_s1.address
		fifo_wrapper_0_s1_write                      : in  std_logic                     := '0';             --                           .write
		fifo_wrapper_0_s1_writedata                  : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		fifo_wrapper_0_s1_read                       : in  std_logic                     := '0';             --                           .read
		fifo_wrapper_0_s1_readdata                   : out std_logic_vector(31 downto 0);                    --                           .readdata
		reset_reset_n                                : in  std_logic                     := '0'              --                      reset.reset_n
	);
end entity fifo_wrapper;

architecture rtl of fifo_wrapper is
	component wrapper is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			avs_s1_address   : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			avs_s1_write     : in  std_logic                     := 'X';             -- write
			avs_s1_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s1_read      : in  std_logic                     := 'X';             -- read
			avs_s1_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			external_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- writebyteenable_n
			external_out     : out std_logic_vector(3 downto 0);                     -- readdata
			ast_source_data  : out std_logic_vector(31 downto 0);                    -- data
			ast_source_error : out std_logic_vector(1 downto 0);                     -- error
			ast_source_valid : out std_logic;                                        -- valid
			ast_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_sink_valid   : in  std_logic                     := 'X'              -- valid
		);
	end component wrapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal fifo_wrapper_0_avalon_streaming_source_valid : std_logic;                     -- fifo_wrapper_0:ast_source_valid -> fifo_wrapper_0:ast_sink_valid
	signal fifo_wrapper_0_avalon_streaming_source_data  : std_logic_vector(31 downto 0); -- fifo_wrapper_0:ast_source_data -> fifo_wrapper_0:ast_sink_data
	signal fifo_wrapper_0_avalon_streaming_source_error : std_logic_vector(1 downto 0);  -- fifo_wrapper_0:ast_source_error -> fifo_wrapper_0:ast_sink_error
	signal rst_controller_reset_out_reset               : std_logic;                     -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal reset_reset_n_ports_inv                      : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv     : std_logic;                     -- rst_controller_reset_out_reset:inv -> fifo_wrapper_0:reset_n

begin

	fifo_wrapper_0 : component wrapper
		port map (
			clk              => clk_clk,                                      --                   clock.clk
			reset_n          => rst_controller_reset_out_reset_ports_inv,     --                   reset.reset_n
			avs_s1_address   => fifo_wrapper_0_s1_address,                    --                      s1.address
			avs_s1_write     => fifo_wrapper_0_s1_write,                      --                        .write
			avs_s1_writedata => fifo_wrapper_0_s1_writedata,                  --                        .writedata
			avs_s1_read      => fifo_wrapper_0_s1_read,                       --                        .read
			avs_s1_readdata  => fifo_wrapper_0_s1_readdata,                   --                        .readdata
			external_in      => fifo_wrapper_0_conduit_end_writebyteenable_n, --             conduit_end.writebyteenable_n
			external_out     => fifo_wrapper_0_conduit_end_readdata,          --                        .readdata
			ast_source_data  => fifo_wrapper_0_avalon_streaming_source_data,  -- avalon_streaming_source.data
			ast_source_error => fifo_wrapper_0_avalon_streaming_source_error, --                        .error
			ast_source_valid => fifo_wrapper_0_avalon_streaming_source_valid, --                        .valid
			ast_sink_data    => fifo_wrapper_0_avalon_streaming_source_data,  --   avalon_streaming_sink.data
			ast_sink_error   => fifo_wrapper_0_avalon_streaming_source_error, --                        .error
			ast_sink_valid   => fifo_wrapper_0_avalon_streaming_source_valid  --                        .valid
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of fifo_wrapper
